module execute(
  input clk_i,
  input reset_i,
  
  input rs1
