module execute(
  input clk_i,
  input reset_i,
  
  input rs1_i,
  input rs2_i,
  input rd_i,
  input aluop_i,
  input 
