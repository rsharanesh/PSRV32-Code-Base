module execute(
