module memory_writeback_register (
    input clk_i, //clock input
    input reset_i, //reset input

    
);
