module memory( 
    input clk_i,//clock input
    input reset_i,//reset input

    
)