module memory_writeback_register (

);
